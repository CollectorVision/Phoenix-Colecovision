--------------------------------------------------------------------------------
--
-- SEX 7264 "COURTNEY"
-- AY-3-8913-COMPATIBLE WSG
-- COPYRIGHT (C) 2019 SILICON SEX
-- HARDCODED BY MADONNA MARK III
--
-- WIP: NATIVE MODE STILL NOT IMPLEMENTED
-- WIP: LEGACY MODE PROVISIONALLY BASED ON THE VERILOG YM2149 CORE WHICH IS
-- COPYRIGHT (C) MIKEJ - JAN 2005
-- COPYRIGHT (C) 2016-2019 SORGELIG
--
-- RELEASED UNDER THE 3-CLAUSE BSD LICENSE:
--
-- REDISTRIBUTION AND USE IN SOURCE AND BINARY FORMS, WITH OR WITHOUT
-- MODIFICATION, ARE PERMITTED PROVIDED THAT THE FOLLOWING CONDITIONS ARE MET:
--
-- 1. REDISTRIBUTIONS OF SOURCE CODE MUST RETAIN THE ABOVE COPYRIGHT NOTICE,
--    THIS LIST OF CONDITIONS AND THE FOLLOWING DISCLAIMER.
--
-- 2. REDISTRIBUTIONS IN BINARY FORM MUST REPRODUCE THE ABOVE COPYRIGHT NOTICE,
--    THIS LIST OF CONDITIONS AND THE FOLLOWING DISCLAIMER IN THE DOCUMENTATION
--    AND/OR OTHER MATERIALS PROVIDED WITH THE DISTRIBUTION.
--
-- 3. NEITHER THE NAME OF THE COPYRIGHT HOLDER NOR THE NAMES OF ITS CONTRIBUTORS
--    MAY BE USED TO ENDORSE OR PROMOTE PRODUCTS DERIVED FROM THIS SOFTWARE
--    WITHOUT SPECIFIC PRIOR WRITTEN PERMISSION.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
--------------------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SEX7264 IS
	PORT
	(
--		 GND															--  1
		 BDIR			: IN  STD_LOGIC						 ;	--  2
		 BC1			: IN  STD_LOGIC						 ;	--	 3
		 DAI			: IN  STD_LOGIC_VECTOR(7 DOWNTO 0); --  4-11
		 DAO			: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --  4-11
--		 TEST_OUT													-- 12
--		 VCC															-- 13
--		 TEST_IN														-- 14
		 DIGITAL_B	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);	-- 15
--		 NO_CONNECT													-- 16
		 DIGITAL_A	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); -- 17
		 DIGITAL_C	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); -- 18
--		 GND															-- 19
		 CLK			: IN  STD_LOGIC						 ;	-- 20
		 CLKENA		: IN  STD_LOGIC						 ;	-- 20*
		nRESET      : IN  STD_LOGIC := '1'            ; -- 21 ON-CHIP PULL-UP
		nA9			: IN  STD_LOGIC := '0'				 ;	-- 22 ON-CHIP PULL-DOWN
		 A8			: IN  STD_LOGIC := '1'				 ;	-- 23 ON-CHIP PULL-UP
		nCHIP_SELECT: IN  STD_LOGIC := '0'				 ;	-- 24 ON-CHIP PULL-DOWN

		 NATIVE		: IN  STD_LOGIC := '0'				 ;	-- 0: LEGACY | 1: NATIVE
--		                                                   (ON-CHIP PULL-DOWN)
		 DIGITAL_MIX: OUT UNSIGNED        (7 DOWNTO 0)	-- MIXED AUDIO
	);
END;

ARCHITECTURE RTL OF SEX7264 IS

-- TYPES

	TYPE PERARRAY  IS ARRAY (1 TO  3) OF STD_LOGIC_VECTOR(11 DOWNTO 0);
	TYPE AMPNARRAY IS ARRAY (0 TO 31) OF UNSIGNED        ( 7 DOWNTO 0);
	TYPE AMPLARRAY IS ARRAY (0 TO 15) OF UNSIGNED        ( 7 DOWNTO 0);

--	CONSTANTS

	CONSTANT AMPLROM : AMPLARRAY :=
	(
		X"00", X"03", X"04", X"06",
		X"0A", X"0F", X"15", X"22", 
		X"28", X"41", X"5B", X"72", 
		X"90", X"B5", X"D7", X"FF" 
	);

	CONSTANT AMPNROM : AMPNARRAY :=
	(
		X"00", X"01", X"01", X"02", X"02", X"03", X"03", X"04",
		X"06", X"07", X"09", X"0A", X"0C", X"0E", X"11", X"13",
		X"17", X"1B", X"20", X"25", X"2C", X"35", X"3E", X"47",
		X"54", X"66", X"77", X"88", X"A1", X"C0", X"E0", X"FF"
	);    

--	SIGNALS

	SIGNAL A			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL B			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL C			: STD_LOGIC_VECTOR(4 DOWNTO 0);

	SIGNAL BC2		: STD_LOGIC := '1'; -- PULLED HIGH INTERNALLY

	SIGNAL BUSADR	: STD_LOGIC;
	SIGNAL BUSENAR	: STD_LOGIC;
	SIGNAL BUSENAW	: STD_LOGIC;

	SIGNAL CLKDIVN	: STD_LOGIC := '0';
	SIGNAL CLKDIVT	: UNSIGNED(3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL CLKENAN	: STD_LOGIC;
	SIGNAL CLKENAT	: STD_LOGIC;

--	TONE DCO'S

	SIGNAL DCOTCNT	: PERARRAY := (OTHERS => (OTHERS => '0'));
	SIGNAL DCOTOUT	: STD_LOGIC_VECTOR( 3 DOWNTO 1) := "000";

--	NOISE DCO

	SIGNAL DCONCNT	: UNSIGNED(7 DOWNTO 0);
	SIGNAL DCONDAT	: STD_LOGIC_VECTOR(16 DOWNTO 0) := (OTHERS => '0');
	SIGNAL DCONOUT	: STD_LOGIC;

	SIGNAL ENVSET	: STD_LOGIC;
	SIGNAL ENVAMP	: STD_LOGIC_VECTOR( 4 DOWNTO 0);
	SIGNAL ENVCNT	: STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL ENVENA	: STD_LOGIC;
	SIGNAL ENVHLD	: STD_LOGIC;
	SIGNAL ENVINC	: STD_LOGIC;
	SIGNAL ENVRES	: STD_LOGIC;

--	INTERNAL REGISTERS

	SIGNAL DCOAPER	: STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL DCOBPER	: STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL DCOCPER	: STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL DCONPER	: STD_LOGIC_VECTOR( 7 DOWNTO 0);

	SIGNAL DCOENA  : STD_LOGIC_VECTOR( 7 DOWNTO 0);

	SIGNAL DCOAAMP : STD_LOGIC_VECTOR( 4 DOWNTO 0);
	SIGNAL DCOBAMP : STD_LOGIC_VECTOR( 4 DOWNTO 0);
	SIGNAL DCOCAMP : STD_LOGIC_VECTOR( 4 DOWNTO 0);

	SIGNAL ENVPER  : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL ENVSHAPE: STD_LOGIC_VECTOR( 3 DOWNTO 0);

	SIGNAL REGADR	: STD_LOGIC_VECTOR( 7 DOWNTO 0);

--	ALIASES

	ALIAS CONTINUE  : STD_LOGIC IS ENVSHAPE(3);
	ALIAS ATTACK    : STD_LOGIC IS ENVSHAPE(2);
	ALIAS ALTERNATE : STD_LOGIC IS ENVSHAPE(1);
	ALIAS HOLD      : STD_LOGIC IS ENVSHAPE(0);

BEGIN

-- BUS CONTROL

-- BDIR BC2 BC1 MODE
-- ---- --- --- -------------
--   0   0   0  INACTIVE
--   0   0   1  LATCH ADDRESS
--*  0   1   0  INACTIVE
--*  0   1   1  READ FROM PSG
--   1   0   0  LATCH ADDRESS
--   1   0   1  INACTIVE
--*  1   1   0  WRITE TO PSG
--*  1   1   1  LATCH ADDRESS

	PROCESS (BDIR, BC1, BC2, A8, nA9, REGADR)
		VARIABLE CS  : STD_LOGIC                   ;
		VARIABLE SEL : STD_LOGIC_VECTOR(2 DOWNTO 0);
	BEGIN
		BUSADR  <= '0';
		BUSENAR <= '0';
		BUSENAW <= '0';

		IF nA9 = '0' AND A8 = '1' AND REGADR(7 DOWNTO 4) = "0000" THEN
			CS := '1';
		ELSE
			CS := '0';
		END IF;

		SEL := BDIR & BC2 & BC1;

		CASE SEL IS
			WHEN "001"	=> BUSADR  <= '1';
			WHEN "011"	=> BUSENAR <= CS ;
			WHEN "100"	=> BUSADR  <= '1';
			WHEN "110"	=> BUSENAW <= CS ;
			WHEN "111"	=> BUSADR  <= '1';
			WHEN OTHERS => NULL          ;
		END CASE;
	END PROCESS;

-- LATCH ADDRESS

	PROCESS (nRESET, BUSADR)
	BEGIN
		IF nRESET = '0' THEN
			REGADR <= (OTHERS => '0');
		ELSIF FALLING_EDGE(BUSADR) THEN
			REGADR <= DAI;
		END IF;
	END PROCESS;

-- LATCH REGISTER

	PROCESS (nRESET, BUSENAW, REGADR)
	BEGIN
		IF nRESET = '0' THEN
			DCOAPER  <=     "111111111111";
			DCOBPER  <=     "111111111111";
			DCOCPER  <=     "111111111111";
			DCONPER  <=         "00000000";
			DCOENA   <=         "11111111";
			DCOAAMP  <=            "11111";
			DCOBAMP  <=            "11111";
			DCOCAMP  <=            "11111";
			ENVPER   <= "1111111111111111";
			ENVSHAPE <=             "1111";
			ENVRES   <=                '0';
		ELSIF FALLING_EDGE(BUSENAW) THEN
			IF NATIVE = '0' THEN
				CASE REGADR(3 DOWNTO 0) IS
					WHEN X"0"   => DCOAPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"1"   => DCOAPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"2"   => DCOBPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"3"   => DCOBPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"4"   => DCOCPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"5"   => DCOCPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"6"   => DCONPER               <= "000" & DAI(4 DOWNTO 0);
					WHEN X"7"   => DCOENA                <= DAI            ;
					WHEN X"8"   => DCOAAMP               <= DAI(4 DOWNTO 0);
					WHEN X"9"   => DCOBAMP               <= DAI(4 DOWNTO 0);
					WHEN X"A"   => DCOCAMP               <= DAI(4 DOWNTO 0);
					WHEN X"B"   => ENVPER  ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"C"   => ENVPER  (15 DOWNTO 8) <= DAI            ;
					WHEN X"D"   => ENVSHAPE              <= DAI(3 DOWNTO 0);
								   ENVRES                <= NOT ENVSET     ;
					WHEN OTHERS => NULL;
				END CASE;
			ELSE
				CASE REGADR(3 DOWNTO 0) IS
					WHEN X"0"   => DCOAPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"1"   => DCOAPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"2"   => DCOBPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"3"   => DCOBPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"4"   => DCOCPER ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"5"   => DCOCPER (11 DOWNTO 8) <= DAI(3 DOWNTO 0);
					WHEN X"6"   => DCONPER               <= DAI(7 DOWNTO 0);
					WHEN X"7"   => DCOENA                <= DAI            ;
					WHEN X"8"   => DCOAAMP               <= DAI(4 DOWNTO 0);
					WHEN X"9"   => DCOBAMP               <= DAI(4 DOWNTO 0);
					WHEN X"A"   => DCOCAMP               <= DAI(4 DOWNTO 0);
					WHEN X"B"   => ENVPER  ( 7 DOWNTO 0) <= DAI            ;
					WHEN X"C"   => ENVPER  (15 DOWNTO 8) <= DAI            ;
					WHEN X"D"   => ENVSHAPE              <= DAI(3 DOWNTO 0);
					               ENVRES                <= NOT ENVSET     ;
					WHEN OTHERS => NULL;
				END CASE;
			END IF;
		END IF;
	END PROCESS;

-- READ REGISTER

	PROCESS (BUSENAR, REGADR , DCOAPER, DCOBPER, DCOCPER , DCONPER, DCOENA,
	         DCOAAMP, DCOBAMP, DCOCAMP, ENVPER , ENVSHAPE)
	BEGIN
		DAO <= "00000000";

		IF BUSENAR = '1' THEN
			CASE REGADR(3 DOWNTO 0) IS
				WHEN X"0"   => DAO <=          DCOAPER ( 7 DOWNTO 0);
				WHEN X"1"   => DAO <= "0000" & DCOAPER (11 DOWNTO 8);
				WHEN X"2"   => DAO <=          DCOBPER ( 7 DOWNTO 0);
				WHEN X"3"   => DAO <= "0000" & DCOBPER (11 DOWNTO 8);
				WHEN X"4"   => DAO <=          DCOCPER ( 7 DOWNTO 0);
				WHEN X"5"   => DAO <= "0000" & DCOCPER (11 DOWNTO 8);
				WHEN X"6"   => DAO <=          DCONPER              ;
				WHEN X"7"   => DAO <=          DCOENA               ;
				WHEN X"8"   => DAO <= "000"  & DCOAAMP              ;
				WHEN X"9"   => DAO <= "000"  & DCOBAMP              ;
				WHEN X"A"   => DAO <= "000"  & DCOCAMP              ;
				WHEN X"B"   => DAO <=          ENVPER  ( 7 DOWNTO 0);
				WHEN X"C"   => DAO <=          ENVPER  (15 DOWNTO 8);
				WHEN X"D"   => DAO <= "0000" & ENVSHAPE             ;
				WHEN OTHERS => NULL                                 ;
			END CASE;
		END IF;
	END PROCESS;

-- CLOCK ENABLE DIVIDERS

	PROCESS (CLK, CLKENA)
	BEGIN
		IF RISING_EDGE(CLK) AND CLKENA = '1' THEN
			CLKENAT <= '0';
			CLKENAN <= '0';

			IF CLKDIVT = "0000" THEN
				CLKDIVT <= "1111";
				CLKENAT <= '1';
				CLKDIVN <= NOT CLKDIVN;

				IF CLKDIVN = '1' THEN
					CLKENAN <= '1';
				END IF;
			ELSE
				CLKDIVT <= CLKDIVT - "1";
			END IF;
		END IF;
	END PROCESS;  

--	NOISE DCO

	PROCESS (CLK)
		VARIABLE DCONCMP  : UNSIGNED(7 DOWNTO 0);
		VARIABLE DCONDAT0 : STD_LOGIC           ;
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF DCONPER  = "00000000" THEN
				DCONCMP := "00000000";
			ELSE
				DCONCMP := UNSIGNED(DCONPER) - 1;
			END IF;

			IF DCONDAT = "00000000000000000" THEN
				DCONDAT0 := '1'; 
			ELSE
				DCONDAT0 := '0';
			END IF;

			IF CLKENA = '1' THEN
				IF CLKENAN = '1' THEN
					IF DCONCNT >= DCONCMP THEN
						DCONCNT <= "00000000";
						DCONDAT <= (DCONDAT(0) XOR DCONDAT(2) XOR DCONDAT0)
						        &   DCONDAT(16 DOWNTO 1);
					ELSE
						DCONCNT <= DCONCNT + 1;
					END IF;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	DCONOUT <= DCONDAT(0);

--	TONE DCO

	PROCESS (CLK)
		VARIABLE DCOTPER : PERARRAY;
		VARIABLE DCOTCMP : PERARRAY;
	BEGIN
		IF RISING_EDGE(CLK) THEN

			DCOTPER(1) := DCOAPER;
			DCOTPER(2) := DCOBPER;
			DCOTPER(3) := DCOCPER;

			FOR I IN 1 TO 3 LOOP
				IF DCOTPER(I)  = X"000" THEN
					DCOTCMP(I) := X"000";
				ELSE
					DCOTCMP(I) := STD_LOGIC_VECTOR(UNSIGNED(DCOTPER(I)) - 1);
				END IF;
			END LOOP;

			IF CLKENA = '1' THEN
				FOR I IN 1 TO 3 LOOP
					IF CLKENAT = '1' THEN
						IF DCOTCNT(I) >= DCOTCMP(I) THEN
							DCOTCNT(I) <= X"000";
							DCOTOUT(I) <= NOT DCOTOUT(I);
						ELSE
							DCOTCNT(I) <= STD_LOGIC_VECTOR(UNSIGNED(DCOTCNT(I)) + 1);
						END IF;
					END IF;
				END LOOP;
			END IF;
		END IF;
	END PROCESS;

--	ENVELOPE FREQUENCY

	PROCESS (CLK)
		VARIABLE ENVCMP : STD_LOGIC_VECTOR(15 DOWNTO 0);
	BEGIN
		IF RISING_EDGE(CLK) THEN
	
			IF ENVPER  = X"0000" THEN
				ENVCMP := X"0000";
			ELSE
				ENVCMP := STD_LOGIC_VECTOR(UNSIGNED(ENVPER) - 1);
			END IF;

			IF CLKENA = '1' THEN
				ENVENA <= '0';
				IF CLKENAT = '1' THEN
					IF ENVCNT >= ENVCMP THEN
						ENVCNT <= X"0000";
						ENVENA <= '1';
					ELSE
						ENVCNT <= STD_LOGIC_VECTOR(UNSIGNED(ENVCNT) + 1);
					END IF;
				END IF;
			END IF;
		END IF;
	END PROCESS;

--	ENVELOPE SHAPE

--     A
-- C   L
-- O   T
-- N A E
-- T T R
-- I T N H
-- N A A O
-- U C T L
-- E K E D
-- -------------
-- 0 0 X X  \___
-- 0 1 X X  /___
-- 1 0 0 0  \\\\
-- 1 0 0 1  \___
-- 1 0 1 0  \/\/
-- 1 0 1 1  \"""
-- 1 1 0 0  ////
-- 1 1 0 1  /"""
-- 1 1 1 0  /\/\
-- 1 1 1 1  /___

	PROCESS (CLK, nRESET)
		VARIABLE ENVBOT  : BOOLEAN;
		VARIABLE ENVBOTP : BOOLEAN;
		VARIABLE ENVTOP  : BOOLEAN;
		VARIABLE ENVTOPM : BOOLEAN;
	BEGIN
		IF nRESET = '0' THEN
			ENVSET <= '0';
		ELSIF RISING_EDGE(CLK) THEN
			IF ENVRES /= ENVSET THEN
				IF ATTACK = '0' THEN
					ENVAMP <= "11111";
					ENVINC <= '0'    ;
				ELSE
					ENVAMP <= "00000";
					ENVINC <= '1'    ;
				END IF;
				ENVHLD <= '0';
			ELSE
				ENVBOT  := (ENVAMP = "00000");
				ENVBOTP := (ENVAMP = "00001");
				ENVTOPM := (ENVAMP = "11110");
				ENVTOP  := (ENVAMP = "11111");

				IF CLKENA = '1' THEN
					IF ENVENA = '1' THEN
						IF ENVHLD = '0' THEN
							IF ENVINC = '1' THEN
								ENVAMP <= STD_LOGIC_VECTOR(UNSIGNED(ENVAMP) + "00001");
							ELSE
								ENVAMP <= STD_LOGIC_VECTOR(UNSIGNED(ENVAMP) + "11111");
							END IF;
						END IF;

						IF CONTINUE = '0' THEN
							IF ENVINC = '0' THEN
								IF ENVBOTP THEN
									ENVHLD <= '1'; 
								END IF;
							ELSE
								IF ENVTOP THEN
									ENVHLD <= '1';
								END IF;
							END IF;
						ELSE
							IF HOLD = '1' THEN
								IF ENVINC = '0' THEN
									IF ALTERNATE = '1' THEN
										IF ENVBOT THEN
											ENVHLD <= '1';
										END IF;
									ELSE
										IF ENVBOTP THEN
											ENVHLD <= '1';
										END IF;
									END IF;
								ELSE
									IF ALTERNATE = '1' THEN
										IF ENVTOP THEN
											ENVHLD <= '1';
										END IF;
									ELSE
										IF ENVTOPM THEN
											ENVHLD <= '1'; 
										END IF;
									END IF;
								END IF;

							ELSIF ALTERNATE = '1' THEN
								IF ENVINC = '0' THEN
									IF ENVBOTP THEN 
										ENVHLD <= '1';
									END IF;

									IF ENVBOT THEN
										ENVHLD <= '0';
										ENVINC <= '1';
									END IF;
								ELSE
									IF ENVTOPM THEN
										ENVHLD <= '1';
									END IF;

									IF ENVTOP THEN
										ENVHLD <= '0';
										ENVINC <= '0';
									END IF;
								END IF;
							END IF;
						END IF;
					END IF;
				END IF;
			END IF;
			ENVSET <= ENVRES;
		END IF;
	END PROCESS;

--	MIX DCOT & DCON

	PROCESS (CLK)
		VARIABLE DCOMIX : STD_LOGIC_VECTOR(2 DOWNTO 0);
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF CLKENA = '1' THEN
				DCOMIX(0) := (DCOENA(0) OR DCOTOUT(1)) AND (DCOENA(3) OR DCONOUT);
				DCOMIX(1) := (DCOENA(1) OR DCOTOUT(2)) AND (DCOENA(4) OR DCONOUT);
				DCOMIX(2) := (DCOENA(2) OR DCOTOUT(3)) AND (DCOENA(5) OR DCONOUT);

				A <= "00000";
				B <= "00000";
				C <= "00000";

				IF DCOMIX(0) = '1' THEN
					IF DCOAAMP(4) = '0' THEN
						A <= DCOAAMP(3 DOWNTO 0) & "1";
					ELSE
						A <= ENVAMP (4 DOWNTO 0);
					END IF;
				END IF;

				IF DCOMIX(1) = '1' THEN
					IF DCOBAMP(4) = '0' THEN
						B <= DCOBAMP(3 DOWNTO 0) & "1";
					ELSE
						B <= ENVAMP (4 DOWNTO 0);
					END IF;
				END IF;

				IF DCOMIX(2) = '1' THEN
					IF DCOCAMP(4) = '0' THEN
						C <= DCOCAMP(3 DOWNTO 0) & "1";
					ELSE
						C <= ENVAMP (4 DOWNTO 0);
					END IF;
				END IF;
			END IF;
		END IF;    
	END PROCESS;

--	MIX CHANNELS

	PROCESS (CLK)
		VARIABLE AUDMIX : UNSIGNED(9 DOWNTO 0);
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF nRESET = '0' THEN
				DIGITAL_A	<= X"00";
				DIGITAL_B	<= X"00";
				DIGITAL_C	<= X"00";
				DIGITAL_MIX	<= X"00";
			ELSE
				IF NATIVE = '1' THEN
					DIGITAL_A <= STD_LOGIC_VECTOR(AMPNROM(TO_INTEGER(UNSIGNED(A))));
					DIGITAL_B <= STD_LOGIC_VECTOR(AMPNROM(TO_INTEGER(UNSIGNED(B))));
					DIGITAL_C <= STD_LOGIC_VECTOR(AMPNROM(TO_INTEGER(UNSIGNED(C))));

					AUDMIX := ("00" & AMPNROM(TO_INTEGER(UNSIGNED(A))))
					       +  ("00" & AMPNROM(TO_INTEGER(UNSIGNED(B))))
					       +  ("00" & AMPNROM(TO_INTEGER(UNSIGNED(C))));

					DIGITAL_MIX	<= AUDMIX(9 DOWNTO 2);
				ELSE
					DIGITAL_A <= STD_LOGIC_VECTOR(AMPLROM(TO_INTEGER(
					             UNSIGNED(A(4 DOWNTO 1)))));
					DIGITAL_B <= STD_LOGIC_VECTOR(AMPLROM(TO_INTEGER(
					             UNSIGNED(B(4 DOWNTO 1)))));
					DIGITAL_C <= STD_LOGIC_VECTOR(AMPLROM(TO_INTEGER(
					             UNSIGNED(C(4 DOWNTO 1)))));

					AUDMIX := ("00" & AMPLROM(TO_INTEGER(UNSIGNED(A(4 DOWNTO 1)))))
					       +  ("00" & AMPLROM(TO_INTEGER(UNSIGNED(B(4 DOWNTO 1)))))
					       +  ("00" & AMPLROM(TO_INTEGER(UNSIGNED(C(4 DOWNTO 1)))));

					DIGITAL_MIX	<= AUDMIX(9 DOWNTO 2);
				END IF;
			END IF;
		END IF;
	END PROCESS;

END ARCHITECTURE RTL;
