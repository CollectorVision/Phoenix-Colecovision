-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity loaderrom is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of loaderrom is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFF5FFFFFFFFFFFFFFFFFFFFFF5FFF5FFF5FFF5FFF5FFF5FFF5F0E7";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4D9F7D";
    attribute INIT_02 of inst : label is "9D4F800D2470B76F4F00036074336001B360F4F5D5B935977649E25CD55B9352";
    attribute INIT_03 of inst : label is "7759D455716B8208D7D532A26E26EEA26A454CA89B89BBAA9A918D774955D776";
    attribute INIT_04 of inst : label is "75498D71D77597B9155655649706D1592511545504565544A28A07860715D767";
    attribute INIT_05 of inst : label is "5494164D5355754D83182733BBEE64944553541575498D549545055D53635855";
    attribute INIT_06 of inst : label is "5455F8F562994626199CA25DB354160575C224152516155D54D0D55E557B9342";
    attribute INIT_07 of inst : label is "5494164D5355755987082733BBEEEE4D575458D549589B75DDA5649706D10592";
    attribute INIT_08 of inst : label is "E4B4BA46D191464270CB2E90E47151517551C2241525161575458D57957B9342";
    attribute INIT_09 of inst : label is "838461E89C14782705391C1463D8E458BA465038D19C463D849E0E118F61270C";
    attribute INIT_0A of inst : label is "A000A000000005FFA497934789C14F1E89C144639162E91EEC671187A2705127";
    attribute INIT_0B of inst : label is "B30BE30000BF800090000008000000080080802A000000000190026090B882BB";
    attribute INIT_0C of inst : label is "E2FBE3FF8255800BE008002202002000000000BFE2F28002F2F822FE22BAA2F8";
    attribute INIT_0D of inst : label is "838FE1BFE02FE2FFE3FFF3FFF3000380B2FFF30033FFF3FC3008330830BF82C0";
    attribute INIT_0E of inst : label is "E2FBE3FF8000000000000000000092002302F00BF3E2F3FFF02FF2FFF00032F8";
    attribute INIT_0F of inst : label is "838FE1BFE02FE2FFE3FFF3FFF3000380B2FFF30033FFF3FC3008330830BF82C0";
    attribute INIT_10 of inst : label is "6904BE65C952500000000000000000000302F00BF3E2F3FFF02FF2FFF00032F8";
    attribute INIT_11 of inst : label is "ECBBBD0555E242497824850915E058D3F8A39EE492EB4907496E45D65C2DCB2F";
    attribute INIT_12 of inst : label is "82B32074941F65055171661ACC81D250759081577756482E4D2492452412FEEB";
    attribute INIT_13 of inst : label is "4B4971F675ECE254D77389505CBFFA45D1C5D65558EB32074941D6E078D21489";
    attribute INIT_14 of inst : label is "9789424978A9346E925E2424978A9346E9258EB32074941D670A413A45C28390";
    attribute INIT_15 of inst : label is "6D2B64931D25D67812FFE9377128576DD1B4AD924B39074975B48915C8555224";
    attribute INIT_16 of inst : label is "F06232141A5BE2C6327D41E73115926F8932414122BA8FEABE63B7B75955DB74";
    attribute INIT_17 of inst : label is "05B9E73250164DECB95BCF264D0152CF5B0C6BAE69649E69505FE1049A0B86BE";
    attribute INIT_18 of inst : label is "24E557ECCD850EF05E0A4D6A3CE8E20627CFCBC7C1F54CDCDCDCD40502B241C5";
    attribute INIT_19 of inst : label is "49754964535496414012F92623676B6F79F54964DB5496497549645354964142";
    attribute INIT_1A of inst : label is "09552550639859362985924198591609859041292623676B6F49F54964DB5496";
    attribute INIT_1B of inst : label is "F263EBBB944DEFE894893944141856041CD55795925E695254956ECEBB2AEC6A";
    attribute INIT_1C of inst : label is "254964D4701505354965CD535AA2AAC94905D505914D505906E49555441B937B";
    attribute INIT_1D of inst : label is "4864254D6A17DB5D354D7FF0E49154955E5050524A07ADEA7A5E857D5418E054";
    attribute INIT_1E of inst : label is "04D5052466254D4AA9BAA062E411515355615925D50464254D6A061158564971";
    attribute INIT_1F of inst : label is "3659649754D645354D641105274DF6EDB76CD525965925D535914D53525D5059";
    attribute INIT_20 of inst : label is "C28504561417541FF0D5795925E6951549FC9299C6254D504149D34199CA25DB";
    attribute INIT_21 of inst : label is "86FE0BF8EF8A24852048D28EFC928ACC6FC93918AFC92A6C68BF244561417141";
    attribute INIT_22 of inst : label is "54D641354D490974919349354D46EF9EE9ED9E254D534E4A464D53524D5350BF";
    attribute INIT_23 of inst : label is "615925D505D64D2464254D5E89388508A6EF9BBA6ED9A254541537DB54D7E417";
    attribute INIT_24 of inst : label is "49354D4E354D4A1049062F496B496749634949F4946B49427494E3494A7F2445";
    attribute INIT_25 of inst : label is "E4A464D53524D53509AEEBBAEEA554D3929193495358BDAD9D8D25392919354D";
    attribute INIT_26 of inst : label is "515254D8BDAD9D8D25392919354D49354D466BBAEEBBA955155362F6B6763494";
    attribute INIT_27 of inst : label is "B1A8254154D151B79535554564979A52908E4A5D53518D53509BBE6EE9BB6689";
    attribute INIT_28 of inst : label is "EBBA95534E4A464D254D62F6B6763494E4A464D53524D53538D53529BB3AECAB";
    attribute INIT_29 of inst : label is "3524DE24D53519AEEBBAEEA554554D8BDAD9D8D25392919354D49354D426BBAE";
    attribute INIT_2A of inst : label is "A54D5290BF8EFE2BF86E824D6EF9BBA6ED9A2545415362F6B6763494E4A464D5";
    attribute INIT_2B of inst : label is "425D2464D24D5350864D5353B76EF9BBA6ED9A25454141151B79535554564979";
    attribute INIT_2C of inst : label is "9362F6B676359F54546B5454275454E35454A460BE413A412896ED9A25551553";
    attribute INIT_2D of inst : label is "4919349354D4619354D4288D059D05AD05BD0564E904A9346924225CAF2BDAFE";
    attribute INIT_2E of inst : label is "54D55515925E694A423929754D46354D42182F904E904A25BB6689554554D097";
    attribute INIT_2F of inst : label is "0B180246554559BB3AECABB1A82541504E2860B6ECEBB2AEC6A09505534546DE";
    attribute INIT_30 of inst : label is "414905712FD27925A4959252495489384107491041D27E617A9E97A12C905710";
    attribute INIT_31 of inst : label is "649525CE262BE6E9B662541527DB5D354171052749E6D4455254BF49E4169056";
    attribute INIT_32 of inst : label is "6156495254DEE41A8A4D649A9AAE649505CAF29050BA41579549C72104501E69";
    attribute INIT_33 of inst : label is "525927B907C99C895254173BFB906EEE41EE41F26722505D525934D525926A45";
    attribute INIT_34 of inst : label is "B3B7BB90706E49F6D74D505F11BDAD9D8D2758593549507EB907B904224E76CD";
    attribute INIT_35 of inst : label is "1D24546DE5415495925E69525FA24E1F11A1191181505DDBFFFFEE4937BFB907";
    attribute INIT_36 of inst : label is "097EE7EA7E67A254963B9C29419C227D505E916D505905D505934D5052924414";
    attribute INIT_37 of inst : label is "C99C8941754964D35496491041D05715541483E6D445525E3BCAC1B421554529";
    attribute INIT_38 of inst : label is "D925B2497BBBBB9279B5115417B9FA719D2541455514A425F8F9FAEBBBBBB907";
    attribute INIT_39 of inst : label is "532495BF35924400C2EEE6495255C8F9355E55EE41CE769E67C9505F9253A495";
    attribute INIT_3A of inst : label is "5556494FBB9A53CE6495055554158FAFDCEE4115256EEEEE41C4F925BA497D92";
    attribute INIT_3B of inst : label is "F6EDBC5117C7E649455157B9749BBC5117C525795055714DD4808F455567D5FD";
    attribute INIT_3C of inst : label is "855D76144926C65BF9A75614492256D4DB1BBC7197C7E649CE76955157B86EF5";
    attribute INIT_3D of inst : label is "A69D967249258E4585124965E1F9A729D115EED55D7197F5445585124A9D6D6D";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD1D610425D55F9E7";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01C";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00BFFC";
    attribute INIT_02 of inst : label is "DC03C01B053CF89C7C0003804B03800AF380C7C8AD4E00AC4780437B8FD4E039";
    attribute INIT_03 of inst : label is "BC4DC2F2C3168902AB880171717531353D02005C5C5D4C4C4F40E00C7D500BC5";
    attribute INIT_04 of inst : label is "1D5084EF00C6D74E000CD51CF20FD6073C71EC0E31E02A88612166A166FCAC10";
    attribute INIT_05 of inst : label is "ECCC00C3B0301D5CA4141A19EC311CF1C7B338401D5884C2355E000754213CD0";
    attribute INIT_06 of inst : label is "EC0D0D02D24FC53F94F493C7C1ECCF008D613C7B33780007558C4308D574E001";
    attribute INIT_07 of inst : label is "ECCC00C3B0301D54A4141A1B6C31D38C01D5884C2351920031B51CF20FC950F1";
    attribute INIT_08 of inst : label is "79FC3043E4AC9B84010F0C10793EA10B2B54A13C7B3378001D5184C23574E001";
    attribute INIT_09 of inst : label is "47C793CD01DCF040771E4F0790E079103040887C21A0790E01DD1F1E43804010";
    attribute INIT_0A of inst : label is "5001522BF00008397800E00F101DCB3CD01DC791E440C107C4681E4F34077077";
    attribute INIT_0B of inst : label is "733D33FFF30070090280000C00A000AE801902D5E380B0000379604902EEE177";
    attribute INIT_0C of inst : label is "330C30307C823334F0B7803301E2D0A280A2834C333C32AD330C33033175F30F";
    attribute INIT_0D of inst : label is "71F4337030303300307E002F430001FB430003FFF00C0304300C330C33407300";
    attribute INIT_0E of inst : label is "330C303070000000000003FFF00903AAB32F73FC007F407E02F4030003FFF30C";
    attribute INIT_0F of inst : label is "71F4337030303300307E002F430001FB430003FFF00C0304300C330C33407300";
    attribute INIT_10 of inst : label is "1E107D3C0FB030000000000000000000032F73FC007F407E02F4030003FFF30C";
    attribute INIT_11 of inst : label is "08423A01565001C0DD00400703F40E217790ED3803268400275384138324871F";
    attribute INIT_12 of inst : label is "658030027500108D4040518600C009D004EA6404C455861584184184184D0084";
    attribute INIT_13 of inst : label is "042760014D75D3EC0C474FB134557784A3010520061803002760135134010040";
    attribute INIT_14 of inst : label is "0D4041C0DC0E000DE025001C0DC0E000DE0261803002760138138403842190E0";
    attribute INIT_15 of inst : label is "21087800809D13544155DE02A01C082B108421E0240E102744E84F0367EAA13C";
    attribute INIT_16 of inst : label is "BC41A6CC0BA4F30D2C2B4890A8CC8B93CC243740314F84F94F81C0BC55420AC4";
    attribute INIT_17 of inst : label is "02EB799EE0038888C88D860CC4ACE30BCEF464F5DF5DF1CFB03B0000E38CC64F";
    attribute INIT_18 of inst : label is "10655BDF824E0F61252F3F6792D25BA5310909090948DFF7FFF7F6DE4B5EC0A8";
    attribute INIT_19 of inst : label is "8C1EC0F8C1EC0F8C6801AE2332F2F2F2D41EC0F8C1EC0F8C1EC0F8C1EC0F8C79";
    attribute INIT_1A of inst : label is "287B136018703E030703E030703E020703E0001E2332F2F2F2E41EC0F8C1EC0F";
    attribute INIT_1B of inst : label is "2309DCC4E4C8888CCE44180C4840169C044302B473D1CFB234C5030A0C2830A1";
    attribute INIT_1C of inst : label is "1EC0F801C07B031EC0F407B03B83E32688007B03E207B03E213845800804E222";
    attribute INIT_1D of inst : label is "6C1D1ECCCC0071C71EC8F5347841EC4C0AD01013040340D0340D02BC80021806";
    attribute INIT_1E of inst : label is "007B033C1F1ECCC24C38C011B801C7B33037473D61201C1ECCCC011C0DD1CF50";
    attribute INIT_1F of inst : label is "1F8C1CF1ECCF801ECCF8031202881F07C1F07B03E1073C7B33E007B333C7B03E";
    attribute INIT_20 of inst : label is "A10087037405848534702B473D1CFB334C50DA4F453ECCE8C480A2014F493C7C";
    attribute INIT_21 of inst : label is "C24F093CE74E00401004C30A50D84A44A50DA6ACE50DA4E45394367037445048";
    attribute INIT_22 of inst : label is "EC8F801EC8CF071CF071CF1ECCCE70F70F70F53EC8E101C1C1C7B133C7B33393";
    attribute INIT_23 of inst : label is "37473D612073C73C1C1EC4DE44184C30E030F0C3C30F13EC8C862071EC8F7801";
    attribute INIT_24 of inst : label is "CF1ECCC21EC4C2310C2312C4D2C4D2C4D2C4D41C4C21C4C21C4CE1C4CE543670";
    attribute INIT_25 of inst : label is "1C1C1C7B233C7B3318320C832061D880707071CFB13C4B4B4B4B910707071EC8";
    attribute INIT_26 of inst : label is "B232188C4B4B4B4B910707071EC8CF1ECCC60C8320C8187B2362312D2D2D2C44";
    attribute INIT_27 of inst : label is "C284A1CCD841C70C3B1300ED1CF473D29381C1C7B13387B13380C3C30F0C3C4F";
    attribute INIT_28 of inst : label is "0C81876201C1C1C73EC4F12D2D2D2E441C1C1C7B233C7B33287B13280C2830A0";
    attribute INIT_29 of inst : label is "233C7D3C7B3338320C832061EC8D88C4B4B4B4B110707071EC8CF1ECCCE0C832";
    attribute INIT_2A of inst : label is "3EC8D39093C24F093C274284030F0C3C30F13EC8C062312D2D2D2E441C1C1C7B";
    attribute INIT_2B of inst : label is "01C73C1C73C7B33081C7B13394030F0C3C30F13EC8C44C1C70C3B1300ED1CF47";
    attribute INIT_2C of inst : label is "E1312D2D2D2D41EC8CA1EC8CA1EC8C61EC8C64823788138810F030F13C7B2363";
    attribute INIT_2D of inst : label is "CF071CF1ECCC6071EC4C6CCB23CB23CB23CB23908E308E208E2083D4F13C4F1D";
    attribute INIT_2E of inst : label is "EC4C03B473D1CF4A4E07071EC4CE1EC4CE30CDE208E2083C0C3C4F1EC8D8C071";
    attribute INIT_2F of inst : label is "00440111AEC0CC0C183060C18461CCD20000003030A0C2830A12871361071C30";
    attribute INIT_30 of inst : label is "C8CF235A08A507333CCC7333CCDA4418C4128C3100A231C0F40D034010612B00";
    attribute INIT_31 of inst : label is "1CFB038D3E4C3F0FC3D3EC0E1071C71EC0F31232800C31C7B13822941C8CF231";
    attribute INIT_32 of inst : label is "3751CFB1348D384927881CF996671CFB134F11E1384D8402B54C1C0781F071CF";
    attribute INIT_33 of inst : label is "B13E234E110CF64FB238800034E231138CD384433D53E207B23E007B23E02470";
    attribute INIT_34 of inst : label is "CBC9CB632013841C71C7B33CB34B4B4B4B3071C30ECCD01DCE134E1091061F07";
    attribute INIT_35 of inst : label is "CA2071C30ECCC37473D1CFB2399106B07B07B07B07B03A0D1C47D38800034E21";
    attribute INIT_36 of inst : label is "095F3FF3DF3FD3EC8EB4F4CFCCF093C7B33DE307B33E307B33E207B339E20C48";
    attribute INIT_37 of inst : label is "0CF64F841EC4F8C1EC4F8C310CA22B4AEC0CEC0C30C3B3363B8E63B0E700ED39";
    attribute INIT_38 of inst : label is "4703B1C0E4C4F4E1030C30EC0D8FE3D8FC3EC8DC03B4E4257EFE7EF64C4F4E11";
    attribute INIT_39 of inst : label is "3B1C0E000073D0D14D3131CFB13E0C3E1C0AD5D38063F8F63F0FB034703B1C0E";
    attribute INIT_3A of inst : label is "4235DF840977E8265DFB037AECCCC3C000D384D0DD5313D384400703B1C0E470";
    attribute INIT_3B of inst : label is "DF37C0B7DC080DFF343F574D08C4C0B7DC1E22B8B0379204AA504FD5408FC3DD";
    attribute INIT_3C of inst : label is "C8D12220A5350B4037FE8220A53FD5137C24C0B7DC080DFFFFD7F03F574C9304";
    attribute INIT_3D of inst : label is "BDF6F7F9DF14209C88294E54E277FD33C71ED310D137DC041C7088294F7D7137";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3F04A20163B6F7F";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFF2FFFFFFFFFFFFFFFFFFFFFF2FFF2FFF2FFF2FFF2FFF2FFF2F01B";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00443F";
    attribute INIT_02 of inst : label is "E097CAB09002011000AAA00A00500AA5000A000300230B337FC25753370230B7";
    attribute INIT_03 of inst : label is "33CE08830B25218D7F230323232727232FC8C0C8C8C9C9C8CBF2DF03CE28F33C";
    attribute INIT_04 of inst : label is "32062CC4F03CE2AF38F5202CB3AB80871CF3FCEF081368A8011124112023021B";
    attribute INIT_05 of inst : label is "FCAC03CFF3B732462CB29CBEAE882CB3CFF2B42732422DFD085708CC838B3103";
    attribute INIT_06 of inst : label is "FCED4C030A4F253C94F293CFE3FCAF0931353CFF2B0021CC90E2C7F4212AF383";
    attribute INIT_07 of inst : label is "FCAC03CFF3B732422CB21CBEAE88ABCA7324A2DFD02B907C0F392CB7AB951830";
    attribute INIT_08 of inst : label is "ABAAEF0AAEEABAABA86ABBC2AAA0F384C082393CFF2B002332282CFD082AF383";
    attribute INIT_09 of inst : label is "AEAAA8194110065044AAA82AA902AAAEEF0BFEEAEAEEAA900ABABAAAA402BA86";
    attribute INIT_0A of inst : label is "F002F11550000270BC29F0805411000194112AAAAABBBC2ABEBBAAA0650442AE";
    attribute INIT_0B of inst : label is "33F4B30041EA90900140000C0350000C00918100107F4009F30F909260CEC3FF";
    attribute INIT_0C of inst : label is "D3AEB2BADC693112F3407033001D03514051430EB30FB150B3AED383B03B4384";
    attribute INIT_0D of inst : label is "B2BAB3AAB2BAB3AAB2AFE2AFE3AAA2BEA380030032AEA1EAD2AEB3AEB3AAB1EA";
    attribute INIT_0E of inst : label is "D3AEB2BAD0000000000003003090015553F43007F2F7E2FEA07EA3AAA000338E";
    attribute INIT_0F of inst : label is "B2BAB3AAB2BAB3AAB2AFE2AFE3AAA2BEA380030032AEA1EAD2AEB3AEB3AAB1EA";
    attribute INIT_10 of inst : label is "2F085E3E4FF0B000000000000000000003F43007F2F7E2FEA07EA3AAA000338E";
    attribute INIT_11 of inst : label is "A8EA6B0BFC7891E2DF88E2478B7E257BB329DABC25B7C207C808C2F327FBC020";
    attribute INIT_12 of inst : label is "F1D9307C882E2F1200002BC764C1F220BCEC707133924A0F42342342342BAA8E";
    attribute INIT_13 of inst : label is "87C882E2111723FC2FFC8FF0BB800BC2CE01928FFF1D9B07C882F3388E2388E2";
    attribute INIT_14 of inst : label is "2DE231E2DE3F0A36F087891E2DE3F0A36F08F1D9B07C882F338FC28FC2F9D9F0";
    attribute INIT_15 of inst : label is "3F8FFC29CF21F30E2E002F0A421623C4F8FE3FF0809F0BC87CE48B8B436AA22E";
    attribute INIT_16 of inst : label is "0232C9101F85F2E349080C38CA109317CB410001345FD5F05F3BEB2364A0F13E";
    attribute INIT_17 of inst : label is "02C8F332140311205009453B84F102321C4E35F2CB0C31C7F0B20101C20CA35F";
    attribute INIT_18 of inst : label is "8A3FF22B44E34F520F4F040057C203243D4D4D4D4F53044448484D00AF820095";
    attribute INIT_19 of inst : label is "C23FC2FC23FC2FC2D401C70A50D0D0F0C33FC2FC23FC2FC23FC2FC23FC2FC2DB";
    attribute INIT_1A of inst : label is "8DBF0B70A87BBF0887BBF0987BBF0A87BBF080170A50D0D0F0C33FC2FC23FC2F";
    attribute INIT_1B of inst : label is "8A952E621ED1120EA6E28D380C2B445422C7FC48B2E2CBF0BAA454A3528D4A34";
    attribute INIT_1C of inst : label is "1FC2FC23C8FF0B3FC2FA4FF0B43209B7C200FF0BF08FF0BF099C2F3FE8121444";
    attribute INIT_1D of inst : label is "8A3E3FC2EA08F3CF3FC2E622FC23FC2FF120A0AAA20BEEFBBEEFBBFA3C2D0422";
    attribute INIT_1E of inst : label is "18FF0B3E3E3FC2D8EAAEA08BBC63CFF0BFC48B2E7A0A3C3FC2EA08BFF122CB9E";
    attribute INIT_1F of inst : label is "3F4D2CB3FC2FC23FC2FC2E030AC23F8FE3F8FF0BD04B2CFF0BF08FF0B3CFF0BF";
    attribute INIT_20 of inst : label is "58822FFC4A29E82622FFC48B2E2CBF0BAA608A4F253FC2D780C2B0994F693CFE";
    attribute INIT_21 of inst : label is "2BECAFB27F27A8EA3A8E69EF60886F2EF608A4AEB608A6B25AD822FFC4AA9E82";
    attribute INIT_22 of inst : label is "FC2FC63FC2CF0F3CF0F3CF3FC2EFC8FC8FC8FC3FC2F083C3C3CFF0B3CFF0BBFB";
    attribute INIT_23 of inst : label is "C48B2E7A08F3CF3E3C3FC2D0E28CE69EF548F523D48F43FC2E1708F3FC2D7C63";
    attribute INIT_24 of inst : label is "CF3FC2E73FC2E7E0269550EAD0EAD0EAE0EAC33EAEB3EAEB3EAE73EAE7D822FF";
    attribute INIT_25 of inst : label is "3C3C3CFF0B3CFF0B9D4952549516DC20F0F0F3CFF0B9434343830F0F0F0F3FC2";
    attribute INIT_26 of inst : label is "F0BA5C29434343834F0F0F0F3FC2CF3FC2E75254952545BF0B70A50D0D0E0D3C";
    attribute INIT_27 of inst : label is "28D236E2DC23CF3CFF0BFF622CB8B2EAAA83C3CFF0B9CFF0B9D523D48F523D0F";
    attribute INIT_28 of inst : label is "52545B7083C3C3CF3FC2E50D0D0E0C3C3C3C3CFF0B3CFF0B9CFF0B9D528D4A35";
    attribute INIT_29 of inst : label is "0B3CF23CFF0B9D4952549516FC2DC29434343834F0F0F0F3FC2CF3FC2E752549";
    attribute INIT_2A of inst : label is "2FC2E9AABB27EC9FB27F27C2548F523D48F43FC2E570A50D0D0E0D3C3C3C3CFF";
    attribute INIT_2B of inst : label is "83CF3C3CF3CFF0B8C3CFF0BBD8548F523D48F43FC2E5623CF3CFF0BFF622CB8B";
    attribute INIT_2C of inst : label is "F0A50D0D0E0C33FC2EB3FC2EB3FC2EB3FC2EBEBAD7C2AFC2ACF548F43DBF0B70";
    attribute INIT_2D of inst : label is "CF0F3CF3FC2E30F3FC2E35439B439B439BC39B0E7F0A7F0A7F0A73FC3B0EC3BC";
    attribute INIT_2E of inst : label is "FC2FFD88B2E2CBAAAA0F0F3FC2E73FC2E7AEB5F0ABF0AB3D523D0F6FC2DC20F3";
    attribute INIT_2F of inst : label is "AF40ABD03FC6C9529D4A7529D276E2D9A79E79E54A3528D4A348DB9B708F3CF3";
    attribute INIT_30 of inst : label is "E6CB9BE75120C79B1E6CB9B2E6FAE28F809AC2E026B0B3EEFEEFBBEE38F0BFA2";
    attribute INIT_31 of inst : label is "1C7F1BE23D163D8F63D3FC2F08F3CF3FC2EE030AC63CF3CFF0BD44831E6C79B2";
    attribute INIT_32 of inst : label is "C480C3F2B00ABC261B412CB6258F2CBF0BC3B8F086EBC2FC44AA3C8F23C8F0C3";
    attribute INIT_33 of inst : label is "F1BD16AF0B80FC0FF1BC6EEEEAF1889945ABC2E03F03F18FF1BF28FF1BF298FF";
    attribute INIT_34 of inst : label is "2C2D2D31B019C63CF3CFF1B96B434343837CF3CF3FC6F092E516AF08B8A33F8F";
    attribute INIT_35 of inst : label is "6B08F3CF3FC6FCC8B2E2CBF0B738A340F40F40F40FF0B70BBAEEABC6EEEEAF18";
    attribute INIT_36 of inst : label is "A90C3CC3DC3DC3FC2D84F2CF2CF6D3CFF1B2F08FF1BF08FF1BF08FF1BEF0B80C";
    attribute INIT_37 of inst : label is "80FC0FC23FC2FC23FC2FC2E022B0BFE3FCAC983CF3CFF0B48D2308C230FF629A";
    attribute INIT_38 of inst : label is "4BABD2EAF2266AF08F3CF3FC2D0F43C0F03FC2C3FD8A6AA4333373732266AF0B";
    attribute INIT_39 of inst : label is "BC2EAFEEECB2D248219882CBF0B4097CBFF112ABC603C0F43D0FF0B0BABC2EAF";
    attribute INIT_3A of inst : label is "A09249EC1451742C041D0993FC2C97FBBBABC20F310899ABC2AFCBABD2EAF0BA";
    attribute INIT_3B of inst : label is "F7BDEABDF6ABBE7917D062AEAC266ABDF6830BFED09935352C093A0E5B0BEE08";
    attribute INIT_3C of inst : label is "EAEAA3538122A9AEF9E65353812D46ABDEA66ABDF6ABBE794F53D3D062AE99AA";
    attribute INIT_3D of inst : label is "04D813604D3A75C1D4E0496A05F9E536CF3DABAAEABDF6AA3CF4D4E04B947ABD";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE4AD2F0009D4135";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFF7FFF7FFF7FFF7FFF7FFF7FFF7F2DF";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0CF0DC";
    attribute INIT_02 of inst : label is "301F00051554555555000150555150055150555F0F44030CCD00604CF1F44031";
    attribute INIT_03 of inst : label is "2CC300F2C0370341F3CD30000C040C0000434C00030103000010C30CC3FF32CC";
    attribute INIT_04 of inst : label is "1FC40B4330CC3D4403F1FF1C7F2EB1071C71CC0C0140001410000700071F0F10";
    attribute INIT_05 of inst : label is "CC0C01C7303F1FC80820342544111C71C730300F1FC80B7C3FD403C7F102D2FF";
    attribute INIT_06 of inst : label is "CC0DC072C2C7071C1C70B1C741CC0D832FC31C3303500FC7FC80BDF3FFD44000";
    attribute INIT_07 of inst : label is "CC0E01C7303F1FC00820742544115100F1FCC0B7C3F435CC330F1C7F2E973071";
    attribute INIT_08 of inst : label is "5554554155555545514515505557C00BC3C4C31C3303500F1F030B7CFFD44000";
    attribute INIT_09 of inst : label is "4545515155545455551555055154555455400054515455154155151545505514";
    attribute INIT_0A of inst : label is "0000000000000EFCD00B40055555451515554551555155055455154545555055";
    attribute INIT_0B of inst : label is "0140400000150100000000000000000000000000000000000050010040010011";
    attribute INIT_0C of inst : label is "0155515501AA4001400000000000000000000001405140005055004150140040";
    attribute INIT_0D of inst : label is "4155505541555055415551555155515550400000015550150155515551555015";
    attribute INIT_0E of inst : label is "0155515500000000000000000100000001401000014051555005505550000041";
    attribute INIT_0F of inst : label is "4155505541555055415551555155515550400000015550150155515551555015";
    attribute INIT_10 of inst : label is "3400131EC7303000000000000000000001401000014051555005505550000041";
    attribute INIT_11 of inst : label is "17052C03FF0432D0C04010CB43010C327D0B45100E190000C7D10030ED9641F0";
    attribute INIT_12 of inst : label is "C34B000C7C030F2FC0C0130D2C0031F00C30D3F1CCFD010C0000000000000140";
    attribute INIT_13 of inst : label is "00C7C0301F0631CC0CC8C73037C00D003B00813FFC34B000C7C0300401004010";
    attribute INIT_14 of inst : label is "0C1002D0C10401034030432D0C1040103403C34B000C7C030C41004100C34B40";
    attribute INIT_15 of inst : label is "0340D00B731F30D90F00340300050CC7340D03400FB400C7CC3007434D40001D";
    attribute INIT_16 of inst : label is "2D07470C04F7C0C307C7C4300C0C84DF0307C3C0407CC7C07CF24C2CF7FF31CD";
    attribute INIT_17 of inst : label is "410F4CE0D404CCCC15C1C72EC4C1F003D0F907C1C71C71C73033C00130DC107C";
    attribute INIT_18 of inst : label is "410FFD73FFC33F71333FC7C01DC087087DC5C5C5C77F547474747F0FC7D0C0C5";
    attribute INIT_19 of inst : label is "001CC0D001CC0D00D000B40303C3C3C3C31CC0D001CC0D001CC0D001CC0D00D2";
    attribute INIT_1A of inst : label is "43F303C010B434000B434000B434000B434000040303C3C3C3C31CC0D001CC0D";
    attribute INIT_1B of inst : label is "340134444C0CCCC1009043EC00043D1400BDFCBC71F1C7303D0FC21008402102";
    attribute INIT_1C of inst : label is "2CC0D000C033031CC0DF073030BB1E19000073034007303401100FFFD4044333";
    attribute INIT_1D of inst : label is "C10D0CC0D00071C71CC0E3D09001CC0FF2F03034100310C4310C433CFC080000";
    attribute INIT_1E of inst : label is "0073031D0C0CC0C7904100021001C7303FC3C71F33010E0CC0D00027F0F1C7CC";
    attribute INIT_1F of inst : label is "1D0C1C71CC0D001CC0D00B0003001D0741D0730343071C730340073031C73034";
    attribute INIT_20 of inst : label is "040009FC3D8CCC03D09FCBC71F1C7303D03C02C7071CC0C2C000C001C70B1C74";
    attribute INIT_21 of inst : label is "D04F413D07D04010040104103C00D00903C03C3D03C02D00740F009FC3D4CCC0";
    attribute INIT_22 of inst : label is "CC0D001CC0C7031C7031C71CC0D060760760761CC0C000C0C0C73031C7303413";
    attribute INIT_23 of inst : label is "C3C71F330071C71D0E0CC0CF904010410C207081C20721CC0D0C0071CC0E1001";
    attribute INIT_24 of inst : label is "C71CC0D41CC0D4B0104303D0C3D0C3D0C3D0C31D0D01D0D01D0D01D0D0CF009F";
    attribute INIT_25 of inst : label is "0C0C0C73031C730353200802008FF000303031C7303C0F0F0F0F0F0303031CC0";
    attribute INIT_26 of inst : label is "3034300C0F0F0F0F0F0303031CC0C71CC0D4C802008023F303C0303C3C3C3C3C";
    attribute INIT_27 of inst : label is "84090FD0F001C71C7303FF2F1C7C71F43400C0C730340730343081C207081C87";
    attribute INIT_28 of inst : label is "08023FC000C0C0C71CC0F03C3C3C3C3C0C0C0C73031C73035073035308402100";
    attribute INIT_29 of inst : label is "031C731C730353200802008FCC0F00C0F0F0F0F0F0303031CC0C71CC0D4C8020";
    attribute INIT_2A of inst : label is "1CC0F43413D04F413D07D000C207081C20721CC0D0C0303C3C3C3C3C0C0C0C73";
    attribute INIT_2B of inst : label is "00C71C0C71C7303500C730340FC207081C20721CC0D0D01C71C7303FF2F1C7C7";
    attribute INIT_2C of inst : label is "40303C3C3C3C31CC0D01CC0D01CC0D01CC0D0D0421004100407C20721FF303C0";
    attribute INIT_2D of inst : label is "C7031C71CC0D4031CC0D4C0F430F430F430F430D04010401040101F4D1344D1F";
    attribute INIT_2E of inst : label is "CC0FFCBC71F1C7D0D003031CC0D01CC0D04108401040101F081C87FCC0F00031";
    attribute INIT_2F of inst : label is "00540015FCC0C30840210084090FD0F41041042C2100840210243F43C0071C71";
    attribute INIT_30 of inst : label is "D0C743C30CC0C7431D0C7431D0F09042C04300B010C030D0F10C4310000033C0";
    attribute INIT_31 of inst : label is "1C7303031CF81E0781E1CC0C0071C71CC0EB0003001C71C7303C33031D0C7431";
    attribute INIT_32 of inst : label is "C3F1C7303C051002CD001C72FCB91C73034D1340010000FCBFD00C0300C031C7";
    attribute INIT_33 of inst : label is "30340144010C74C73030044454401111005100431D31C0073034007303400B9F";
    attribute INIT_34 of inst : label is "858585801011001C71C73038300F0F0F0F0C71C71CC0F0134401440124101D07";
    attribute INIT_35 of inst : label is "0C0071C71CC0FC7C71F1C73032E4103C33C33C33C33032C11846510044454401";
    attribute INIT_36 of inst : label is "43DF1DF1DF1DF1CC0D0C70070070F1C73033400730340073034007303F402C00";
    attribute INIT_37 of inst : label is "0C74C7001CC0D001CC0D00B010C033CFCC0C0B1C71C730364190641905FF2F43";
    attribute INIT_38 of inst : label is "4B4352D0D4445440071C71CC0D8761D8761CC0D7FCBD0D0F7D7D7D7D44454401";
    attribute INIT_39 of inst : label is "352D0D444471C000011111C73031C1F027F2FF510061D8761D873034B4352D0D";
    attribute INIT_3A of inst : label is "FFF1C7C80071F0081C7303FFCC0C1F111151005F1FD11151000A8B4352D0D4B4";
    attribute INIT_3B of inst : label is "DD374177DC151DF7D7CBFD47F0044177DC14033C303FF000C400265FFFDFCB5B";
    attribute INIT_3C of inst : label is "57F3FF00010D15F477DF3F00010DFD3F74544177DC151DF76DDB7FCBFD45510F";
    attribute INIT_3D of inst : label is "2C74B1D2C70F1057C00041DF4577DC07871C513FF3F7DC0F1C7FC0004377D3F7";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB01009007FF4B1D";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
